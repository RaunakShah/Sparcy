module top
#(
  BUS_DATA_WIDTH = 64,
  BUS_TAG_WIDTH = 13
)
(
  input  clk,
         reset,

  // 64-bit address of the program entry point
  input  [63:0] entry,
  
  // interface to connect to the bus
  output bus_reqcyc,
  output bus_respack,
  output [BUS_DATA_WIDTH-1:0] bus_req,
  output [BUS_TAG_WIDTH-1:0] bus_reqtag,
  input  bus_respcyc,
  input  bus_reqack,
  input  [BUS_DATA_WIDTH-1:0] bus_resp,
  input  [BUS_TAG_WIDTH-1:0] bus_resptag
);

  // instantiate processor core
  Core #(64, 13) core(
    clk, reset, entry,
    bus_reqcyc, bus_respack, bus_req, bus_reqtag,
    bus_respcyc, bus_reqack, bus_resp, bus_resptag
  );

  initial begin
    $display("Initializing top, entry point = 0x%x", entry);
  end
endmodule
