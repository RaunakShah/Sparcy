`ifndef __alu__ops
`define __alu__ops

// macro definitions for op3 

`define ADD 3'b101 // need to change this one too

`endif

